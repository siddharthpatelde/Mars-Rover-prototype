PK   sW�-U�  ��     cirkitFile.json�]��F��+\-�,Dm?�ds�r@�M6�ǭ�8�!4ɦ��8�(?����p��)J")��qS�A����__UW���'�z���8/���.VY��\R1�\�"y��o�tr�-�e>U�����{���n��7��R/˹�L��f�Va�z�`n��b�P����zN&�/�UN���<fnPY��U�Wn���+�2	������[�6-���M˲�e��$I�K]/P"�':�4f!M�3ۨ��l[T������|?�]���b�s�P�ya��j��	���� ��p�j�j�Yh�4?�J�s���)`,NCWzJB�2`:��"�yVղ�J6M�^�DU?�j�P��q���p�$u#�.p�T�؏�8�*ô|��ղ�X�I%�e�T�Įz�恓��c�zi��3�]�F2m��>�0��+����x��.!D�� _ J,VIج�X%n�J=u�Z��;Z�HqS�Y��ĩ����L(���P�Xab�¾�vե��͸Þ��;��ڶU��z�Z*~j���gY_Xַ�<��<������R4V���.�3Qz�J�%�%�%�%�%�YгtHWΦ�]/�i�O֐���R�x�6���!.O(
?��M�0���|qॱpNP�-[�VT�~aEU�UT�~QEڂg𤑛�E˴?��2b��D9Hg	e�64� (��/q���/�?+B4��]�׃ɟI
��,�0�%M� =.6�?<"l�FT�X��'�t6�nf7��jD�  o+W�ļ`C���7��)-��Sx����>!���}��%�I�m�h���b�#p9��Q���3/�)�`c��x�ƥFQ0
yj?�F��% =�㠗�_:~�71�q L��0�㰩P&�m����bV�8H"a�f�qP��A1�l���u���ΰ��ь�y���؀�\���I��FqF�rR��1�a.��ΰm���`l��O�����Iq����5V�*�mPc��e��A{.�tPÞ�����\�A{.'G�j�s᧸���\N�:�a��传��\NK 6�a��传��\N�:�a�e�y�F�"F���%���K8�F�8������_:��8��@���a:��8(f㠘����A1�l�qP��A1�l�qP��A1?�btPÞ�8}9)P蠆=���jrA5� <8dPÞ�8}i����|[n�4�Y�vrI�t�&+�j~�P�N��r��.&�/i!QNe��"��4M��R��i����B����9o���Z�̹�[=���c�d㜞�ed��-#�`�u���l3f�*�r�����3����a��9ƌ��`��;��k���G{�FF?��O���F�;���M���e��c岞A����YvJ�A�3�n�!J��+Vр�/��b�o��`)�er�h|��{�}�k��^T\,zQ��������`>�A}�`��u k^�c��ʶ�Kc�l���g� ��>���f i�#��Ok�v����=�$ֺ}l���|
�}��Ą?�n�Z�gܢq���]B>�yo|�/��r��{��t�K�[g�m:i�� ��a�c���:�l����N��[&��&�5�:}�����>2X+����Y��;t�]�]�D�\�����p��N�C�6�n���o���3��<��J�wgS�v�,�;X��w6�,�K��N��a��g^[�R[�R[�V�vV�-[�R[�V9uV� 3�M��ҊG6i�Yg�![�2[�2[�2[�V�s�E�1��It~VgB���ǆŧ�Y����JgS߶��A'����t�\O}t�ΚA���,:q�;t]�[��L�;����=�,1�2L��\�d�h�U�Ԇ��*a�v���d|M0��ъO�hE��9�8��gT��.���iqӊ�PRCJ-5��PSCN=5���LV�65���Lfj0S����`�FuW����i��F����=�@H���-1�=x����a����l#��v����K]��7����e�vW�ll��6�� ���j��r�*-��<��6_���r�O�t��[�gm�txhN[��j��xh<[ݤj��x�X])k��x�����.��Њ��^�2���̳�1����~�.�ፅ���lՇ{��.��5yUD�X]��x]�����;,u�8,��"��(����"YU��Z,�\�l���E�*����|>g���Z�A�ڳ4g,��͟�B���CO�/����T��}��i���̴��e"�*+�����,�>�|"|����tF2泀��38�<[�{��>l@I�R"��F^B=����!�:J��7uP��t�t]mz6Y�«8+Ⅾ��e$�y�9����x	'3�!������N�3��`�>��Uÿf�r�d����nBgtF`�L���vi~���UYd�W0���1Ϧt:y�k���#.��X/3X�	�����<Y> ���T-V
W��9[e�B����uVh��pky���T����P�M�}G��j�<��*�77#��0@���'y=߾7��g�/|���FT�����A�4I��0���+'!]`���.����uy�-��� A -^��h������]/��f!�L�&<;��}�إB��g��g������rt`�4 3�'^O�S�X8�����EW$H��C�	�ƮT���,P� `�ֺ�-T�-�A
�wd���'Ϙ�{녂�p3�	�f���$ M5IhH<�Ezp9;���?H}���Xg%�dm���ՖK	�	��{�mb���[�Еʔ'
0E`[wYE���{�)(4�%����j.�:%�T��!�J(i>1Ѳ5�'�?]�I�SIwe���>�R���7!�qfW�
�A�>@�G���2Jb�C��&ʉUH��`��+��'�*�����p��2�?U��9%�3�(�,h-�0�D7���΃",��Û@�ǺAų��e�K�����i��O�4�(m���徴ʶ`:V�xͲz��>�&%�2�*�[eE�Z7�V_d����2�o>���@a=�>gi[�H�'����9K��o�X����D��o���W^�� 4����"����U%�W�˫��W]��W���$K�7<�-4	��D��c 	�X���AE���.r�ʛ��M]0⸦R����E<���������k�oԋS�s/��e��(��)r�T������{��]���R�T���r����&$�J��X�$�1��p�p�OmX<�9����H\g����D�<�㗸����P\��0Hh/�ZS�@E^>����qIp���w�0��6�>�҈K�IM�#\,�n�3�x�)��0Ĉ����Ei�H��woo�2Ѧ�Q��N����1��-ZV+�f��-,jM����I��i^��$I�W����)��'�4[�#ȚA�&���-N���sv���D�£�$��}҇.�4u�j������}�`�*�G�E��|��~BaŮ�<�R�ƚ�A,�E�H��\�� MBc�f��<��i��t]���j��l/։v���?<�]����r��.^�ݗ���m^����L/Wyᘏ̆,�i��0{���9����R'�^e�Z�������a5�O��P�|���wPԡ�]�����ϡ�C��R-�W�j�o�� �wT��C�.`�k�!��<;����CΣ��qiF�s���b3��f�_�JLc7���f?���V�U�)��lYօ_;?>��Ԉs��S��]��_;���Vf��"b��5tn�U��������-�unL���<K[|�g�Gy�2��E��]Q5�λ�"l�S�p�}5�fɶp�����W�{x��|��,f�~�-/B���v���r������<�XGm�̫�.MY-:s̀�툇�٬��s}�25 Q����&K���pu>kbv3��ެ�?�
E.f5t0�����mV6� ��T�/j��TY���b����薋(�Γ��?��y�|+]S���m�ƒ/�|��Y�\ԝU�U�0b���-�S��,�Nj��z7BU�@k��!�]q�=C�z���t)v�:N�Vڡ��g�Gb��&X�����Y�zC����n��7����H�P]ѭ{ �C��f��޺"�[�.����8����J���[�P��.�j�(O���%�ŕ~�h����v�=���^�l9�͆�P��Б�C���J�M[?w|'�G��O��|�<���,j}L�|��k�p���5��t�Fh���U�@7+�S^k�e�h������n�غ��Pl�aoXh����k�o2�"^��x}h��i��xc�_|C�nYU[#��ԺtZm�o;�;�D/ԻJv��11�����uL�6K�E�����(_�"W�s�k�Y��I�/���l�4&�K���U�k��fVK������׿���e����&���{��N��q�"�1]��O��8�^�3 ��鸉ǯK��V��e��^�S�z�T��>ͳ�����U\��41:Ĥ�g���`�b:T�{�1�����!�?���A[-���e�:�І���A&뢊��mg%�&��1��������?/]]G)����*�75Q��=��"_�8_&��/;Z�����a�:%'�Z� x�^�]�!�n;�\���������:�W����7��������Q>'����p����N�O��M�+JѴ�E�|�2����졿8�g����ol���g� �����c��q�(y�d_P�H��y��I=0x�I�)����L�O�����UG�XT#�8���*�4<�i6�E�|�+��^�~���*���ֱ�cַ&���� �B��O]O�e�4>��l���7�{S烣�|n�q����l�i)uo4=�6ߪ�՟\���[d:���h�<�$OI���/>&+���%�?�\�]��ɐ�g�0���P��i�]���%~�R3�2.��O��v��P�u1� �I3�R���2%D����)f<d�o2��PxT�,4B�^
Nf~ �O��3B<���	_�GYe�|t���4��o�M��ҿE �sC�0̱!Y�^����09�ҍ�� �.�f�Z�E� V�uN��t�.�PJ�2t���Yrv���ɷ.��/>���ٌz��b+��f�A^�3����Q��P	�5�]��p�dZ]�9�� ����Y��6����H4�ԙM˱�د>��N�KwJ_�C�>yi9�p4�\ԟ[[x=���|-���{�[�ƛz�1�A)h74����������,�%+���ڮ*Ao"������������w�K��EZ�x_�ɭ��#?�Ȗj�do����}_���F��:͗��w}��p�Gr�[/�F��k���X��^����^�l?�e��Ō�>�@`�-�[��E��0ty��%w}�*���g���ꪒ�j��2�x*EU���#���S�A��	�b
��F��ɒ��pؤwܜ���U�>�fF��g�@��V}�bo�R�N��#~Z�|�s���b�Qs~���8m�DI
8�$�d f�:���4٤�.�AV��F*V�z�l̮�����m*��*�+^�weNm?I���g��T�\�/���c�{�i�<�̈��%�'��d���;�Qp:t/�Y� ��@{A��v���5�}�o���?<p�)�<�е{V�c¢Z���ւv�����yu/�C����=L��؂v���@]kv?��w�7��޲��B�'��,뎻��^��]��uo��̂�.��~Rss��=�����Wq���YO��pd>8�G�!�� l�M����`�Fvl��7�c۳�gvlym#�w齠�]�_tt�P�
g�kρ�]����;t�uo/#=ʃ���J�{���v�������8�_{x�n}�x�v�{Kǯ���ҝi��ܺ}O��k���]��`���78��ݛ�V?li�ac�7#����͸�39�{ӺZ�wݑd�O�t=�"R��ߌ��X0��3�2��g��=&��2s1�Q:���;�a��1]��G�q�U u�>�㝹��x�����~G�t=[�D������z�c�;�1w��h��M���/�^z,?�m r@w"	ORN��G�"wP"w��X�H�����ʎ}����f��6C���oDB;�m,�Џ�H;�~�k_���X"��^c�HHQ�搮Ϥ�H��^�i�лlG辍��Q�t���#�(�Z(��m bRm���I�H�Ձ����`fU=d���Z������a�o�-�/^~�|�?PK
   sW�-U�  ��                   cirkitFile.jsonPK      =       